tb_ace_ccu_top.sv